//`define         PLATFORM_GENERIC          1
`define         PLATFORM_ALTERA           1
//`define         PLATFORM_XILINX           1
`define ZUMA_LUT_SIZE 5