`define         PLATFORM_XILINX           1
