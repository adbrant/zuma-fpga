`define ZUMA_LUT_SIZE 6
